module queue();
// function queue,
// do one thing per cycle.

endmodule
