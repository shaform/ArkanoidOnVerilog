module word(
	input [4:0] row, col,
	input [1:0] select,
	output word
);
reg [19:0] data;
always @(row,col,select,data[19:0])
begin 
	case (select)
		2'b00: case(row) // waiting to start.
				5'b00000: data = 20'b00000000000000000000;
				5'b00001: data = 20'b00000111111111100000;
				5'b00010: data = 20'b00011000000000011000;
				5'b00011: data = 20'b00100000000000000100;
				5'b00100: data = 20'b01000111000011100010;
				5'b00101: data = 20'b01001000100100010010;
				5'b00110: data = 20'b01000000000000000010;
				5'b00111: data = 20'b01000100000000100010;
				5'b01000: data = 20'b00100011111111000100;
				5'b01001: data = 20'b00011000000000011000;
				5'b01010: data = 20'b00000111111111100000;
				5'b01011: data = 20'b00000000000000000000;
				5'b01100: data = 20'b00000000000000000000;
				5'b01101: data = 20'b00011111000011110000;
				5'b01110: data = 20'b00100000000100001000;
				5'b01111: data = 20'b00100000001000000100;
				5'b10000: data = 20'b00100111101000000100;
				5'b10001: data = 20'b00100011000100001000;
				5'b10010: data = 20'b00011110000011110000;
				5'b10011: data = 20'b00000000000000000000;
				default: data = 20'bxxxxxxxxxxxxxxxxxxxx;
			endcase
		2'b01: case(row) // lose
				5'b00000: data = 20'b00000000000000000000;
				5'b00001: data = 20'b00100011101110111000;
				5'b00010: data = 20'b00100010101000100000;
				5'b00011: data = 20'b00100010101110111000;
				5'b00100: data = 20'b00100010100010100000;
				5'b00101: data = 20'b00111011101110111000;
				5'b00110: data = 20'b00000000000000000000;
				5'b00111: data = 20'b00001110000001110000;
				5'b01000: data = 20'b00011111000011111000;
				5'b01001: data = 20'b00011111110001111000;
				5'b01010: data = 20'b00001111100111110000;
				5'b01011: data = 20'b00000011110001100000;
				5'b01100: data = 20'b00000001100001000000;
				5'b01101: data = 20'b00000000100000000000;
				5'b01110: data = 20'b00011110000000000000;
				5'b01111: data = 20'b00100000111100100100;
				5'b10000: data = 20'b00011100100010100100;
				5'b10001: data = 20'b00000010111100011100;
				5'b10010: data = 20'b00000010100010000100;
				5'b10011: data = 20'b00111100100010011000;
				default: data = 20'bxxxxxxxxxxxxxxxxxxxx;
			endcase
		2'b10: case(row) // nothing
				default: data = 20'bxxxxxxxxxxxxxxxxxxxx;
		       endcase
		2'b11: case(row) // win
				5'b00000: data = 20'b00000000000000000000;
				5'b00001: data = 20'b01000001000000000010;
				5'b00010: data = 20'b00101010010011100010;
				5'b00011: data = 20'b00101010000010010010;
				5'b00100: data = 20'b00111110010010010000;
				5'b00101: data = 20'b00010100010010010010;
				5'b00110: data = 20'b00000000000000000000;
				5'b00111: data = 20'b00100010011000001100;
				5'b01000: data = 20'b00010100100100010010;
				5'b01001: data = 20'b00001000100100010010;
				5'b01010: data = 20'b00001000100100010010;
				5'b01011: data = 20'b00001000011001001100;
				5'b01100: data = 20'b00000000000000000000;
				5'b01101: data = 20'b00000000000000000000;
				5'b01110: data = 20'b00000000000000000000;
				5'b01111: data = 20'b00000000000000000000;
				5'b10000: data = 20'b00000000000000000000;
				5'b10001: data = 20'b00000000000000000000;
				5'b10010: data = 20'b00000000000000000000;
				5'b10011: data = 20'b00000000000000000000;


				default: data = 20'bxxxxxxxxxxxxxxxxxxxx;
		       endcase
		default: data = 20'bxxxxxxxxxxxxxxxxxxxx;
	endcase
end

assign word = data[19-col];

endmodule
