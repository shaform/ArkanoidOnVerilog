module block_select(
	input blocks,
	input [6:0] row, col,
	output [3:0] block
);
endmodule
