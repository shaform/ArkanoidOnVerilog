module test_ball(
);

reg [9:0] x, y;


always @(posedge clock)
begin
	if (reset) begin
		x <= 40;
		y <= 80;
		x_ang <= ;
		y_ang <= ;
	end else begin
	end
end




endmodule
