module draw_block(
	input vcounter,
	input hcounter,
	output [3:0] out
);

endmodule
